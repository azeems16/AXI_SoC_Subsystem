class soc_timer_coverage